module nsubburaj_lab1_verilog(a,b,Y);
input a,b;
output Y;
assign Y = a & b;
endmodule