module nsubburaj_lab2_verilog(a,b,Y);
input a,b;
output Y;
assign Y = a | b;
endmodule